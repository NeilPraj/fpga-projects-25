//

module QuadDecoder (
    input logic clk, 
    input logic rst_n, 
    input logic [15:0] bcd_in, 
    output logic [6:0] seg_out, // 7-segment display output
    output logic [3:0] digit_select // Digit select for multiplexing
);
    



endmodule